CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
310 140 8 100 10
241 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
5 4 0.323838 0.500000
409 176 522 273
244318226 0
0
6 Title:
5 Name:
0
0
0
101
13 Logic Switch~
5 112 377 0 10 11
0 113 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5582 0 0
2
42755.5 0
0
9 Inverter~
13 783 333 0 2 22
0 4 3
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U27F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 16 0
1 U
5236 0 0
2
5.89785e-315 0
0
9 Inverter~
13 839 486 0 2 22
0 7 6
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U27E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 16 0
1 U
348 0 0
2
5.89785e-315 0
0
9 2-In AND~
219 834 415 0 3 22
0 4 6 5
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U18A
-37 -25 -9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6515 0 0
2
5.89785e-315 0
0
9 2-In AND~
219 744 436 0 3 22
0 4 7 8
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U29D
-37 -25 -9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
9161 0 0
2
42755.5 1
0
9 2-In XOR~
219 127 198 0 3 22
0 11 10 9
0
0 0 608 180
6 74LS86
-21 -24 21 -16
3 U3D
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6245 0 0
2
42755.5 2
0
9 Inverter~
13 57 198 0 2 22
0 9 12
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U27D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 16 0
1 U
9279 0 0
2
42755.5 3
0
2 +V
167 1454 211 0 1 3
0 19
0
0 0 54240 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5268 0 0
2
42755.5 4
0
5 4073~
219 1238 46 0 4 22
0 15 14 13 20
0
0 0 608 180
4 4073
-7 -24 21 -16
4 U17A
-16 -25 12 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 20 0
1 U
3891 0 0
2
42755.5 5
0
5 4081~
219 1391 72 0 3 22
0 14 13 18
0
0 0 608 180
4 4081
-7 -24 21 -16
4 U19D
-16 -25 12 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
9369 0 0
2
42755.5 6
0
9 Inverter~
13 1293 596 0 2 22
0 25 43
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U4F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
8239 0 0
2
42755.5 7
0
9 Inverter~
13 1325 594 0 2 22
0 25 42
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U27A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
7160 0 0
2
42755.5 8
0
9 Inverter~
13 1261 592 0 2 22
0 25 44
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U27B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 16 0
1 U
9517 0 0
2
42755.5 9
0
9 Inverter~
13 1229 594 0 2 22
0 25 45
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U27C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 16 0
1 U
7689 0 0
2
42755.5 10
0
7 Ground~
168 919 595 0 1 3
0 2
0
0 0 53344 270
0
5 GND13
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3436 0 0
2
42755.5 11
0
2 +V
167 917 572 0 1 3
0 46
0
0 0 54240 90
2 5V
-7 -15 7 -7
3 V16
-10 -25 11 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7951 0 0
2
42755.5 12
0
7 Ground~
168 951 522 0 1 3
0 2
0
0 0 53344 270
0
5 GND14
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3710 0 0
2
42755.5 13
0
9 2-In AND~
219 1192 556 0 3 22
0 30 25 35
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U13B
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3654 0 0
2
42755.5 14
0
9 2-In AND~
219 1096 555 0 3 22
0 33 25 41
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U13C
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
7865 0 0
2
42755.5 15
0
9 2-In AND~
219 1128 555 0 3 22
0 32 25 39
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U13D
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3647 0 0
2
42755.5 16
0
9 2-In AND~
219 1160 556 0 3 22
0 31 25 37
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U28A
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
8917 0 0
2
42755.5 17
0
9 2-In AND~
219 1288 557 0 3 22
0 23 43 36
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U28B
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
9355 0 0
2
42755.5 18
0
9 2-In AND~
219 1256 556 0 3 22
0 22 44 38
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U28C
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
7514 0 0
2
42755.5 19
0
9 2-In AND~
219 1224 556 0 3 22
0 21 45 40
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U28D
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
7418 0 0
2
42755.5 20
0
9 2-In AND~
219 1320 557 0 3 22
0 24 42 34
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U29A
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
4510 0 0
2
42755.5 21
0
8 2-In OR~
219 1141 495 0 3 22
0 41 40 26
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U11B
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5695 0 0
2
42755.5 22
0
8 2-In OR~
219 1176 496 0 3 22
0 39 38 27
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U11C
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
7349 0 0
2
42755.5 23
0
8 2-In OR~
219 1209 497 0 3 22
0 37 36 28
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U11D
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3818 0 0
2
42755.5 24
0
8 2-In OR~
219 1244 498 0 3 22
0 35 34 29
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U30A
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
629 0 0
2
42755.5 25
0
4 4008
219 1005 564 0 14 29
0 2 22 23 24 46 46 46 2 122
30 31 32 33 123
0
0 0 13024 0
4 4008
-14 -60 14 -52
3 U31
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3663 0 0
2
42755.5 26
0
9 2-In AND~
219 933 435 0 3 22
0 21 22 48
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U29C
-37 -25 -9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
9622 0 0
2
42755.5 27
0
9 2-In AND~
219 969 436 0 3 22
0 21 23 47
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U29B
5 -26 33 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
7514 0 0
2
42755.5 28
0
8 2-In OR~
219 947 380 0 3 22
0 48 47 25
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U30B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
5133 0 0
2
42755.5 29
0
7 Pulser~
4 1558 268 0 10 12
0 124 125 49 126 0 1 99 66 22
8
0
0 0 4640 512
0
3 V15
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3505 0 0
2
42755.5 30
0
12 D Flip-Flop~
219 1457 299 0 4 9
0 16 49 127 21
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 Qd
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4860 0 0
2
42755.5 31
0
12 D Flip-Flop~
219 1371 299 0 4 9
0 15 49 128 22
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 Qc
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5298 0 0
2
42755.5 32
0
12 D Flip-Flop~
219 1277 299 0 4 9
0 14 49 129 23
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 Qb
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4443 0 0
2
42755.5 33
0
12 D Flip-Flop~
219 1193 300 0 4 9
0 13 49 130 24
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 Qa
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8393 0 0
2
42755.5 34
0
7 Pulser~
4 1084 85 0 10 12
0 131 132 17 133 0 0 33 22 22
8
0
0 0 4640 0
0
3 V14
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5166 0 0
2
42755.5 35
0
2 +V
167 1121 211 0 1 3
0 19
0
0 0 54240 180
2 5V
7 -2 21 6
3 V13
4 -12 25 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
818 0 0
2
5.89785e-315 0
0
5 4027~
219 1495 184 0 7 32
0 134 19 17 19 135 136 13
0
0 0 4704 0
4 4027
7 -60 35 -52
2 Qa
30 -61 44 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 15 0
1 U
4292 0 0
2
5.89785e-315 5.26354e-315
0
5 4027~
219 1400 184 0 7 32
0 137 13 17 13 138 139 14
0
0 0 4704 0
4 4027
7 -60 35 -52
2 Qb
30 -61 44 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 15 0
1 U
33 0 0
2
5.89785e-315 5.30499e-315
0
5 4027~
219 1301 184 0 7 32
0 140 18 17 18 141 142 15
0
0 0 4704 0
4 4027
7 -60 35 -52
2 Qc
30 -61 44 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 14 0
1 U
9412 0 0
2
5.89785e-315 5.32571e-315
0
5 4027~
219 1193 184 0 7 32
0 143 20 17 20 144 145 16
0
0 0 4704 0
4 4027
7 -60 35 -52
2 Qd
30 -61 44 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 14 0
1 U
3792 0 0
2
5.89785e-315 5.34643e-315
0
7 Ground~
168 754 647 0 1 3
0 2
0
0 0 53344 90
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7568 0 0
2
5.89785e-315 5.3568e-315
0
7 74LS181
132 702 687 0 22 45
0 53 2 2 53 11 52 51 50 21
22 23 24 146 2 4 147 148 149 61
60 59 58
0
0 0 4832 0
6 74F181
-21 -69 21 -61
3 U22
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3380 0 0
2
5.89785e-315 5.36716e-315
0
2 +V
167 647 627 0 1 3
0 53
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V12
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8942 0 0
2
5.89785e-315 5.37752e-315
0
7 Ground~
168 663 627 0 1 3
0 2
0
0 0 53344 180
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4537 0 0
2
5.89785e-315 5.38788e-315
0
6 74LS85
106 819 637 0 14 29
0 54 55 56 57 61 60 59 58 150
151 152 153 7 154
0
0 0 5088 0
5 74F85
-18 -52 17 -44
3 U14
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9868 0 0
2
5.89785e-315 5.39306e-315
0
4 LED~
171 753 243 0 2 2
12 8 2
0
0 0 880 180
4 LED1
-30 7 -2 15
3 WIN
-24 -14 -3 -6
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8516 0 0
2
5.89785e-315 5.39824e-315
0
4 LED~
171 807 243 0 2 2
10 5 2
0
0 0 880 180
4 LED1
8 7 36 15
4 LOSE
6 -14 34 -6
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7565 0 0
2
5.89785e-315 5.40342e-315
0
4 LED~
171 784 273 0 2 2
11 3 2
0
0 0 880 180
4 LED2
6 7 34 15
3 OVF
4 -14 25 -6
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8189 0 0
2
5.89785e-315 5.4086e-315
0
7 Ground~
168 783 204 0 1 3
0 2
0
0 0 53344 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4137 0 0
2
5.89785e-315 5.41378e-315
0
8 Hex Key~
166 672 241 0 11 12
0 57 56 55 54 0 0 0 0 0
15 70
0
0 0 4640 512
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3419 0 0
2
5.89785e-315 5.41896e-315
0
9 CC 7-Seg~
183 928 137 0 17 19
10 77 76 72 71 73 74 75 155 2
0 1 1 0 0 0 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8648 0 0
2
5.89785e-315 5.42414e-315
0
9 CC 7-Seg~
183 1026 138 0 17 19
10 70 69 68 64 65 66 67 156 2
1 0 1 1 0 1 1 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7219 0 0
2
5.89785e-315 5.42933e-315
0
4 4511
219 921 241 0 20 29
0 157 158 159 25 2 63 63 75 74
73 71 72 76 77 0 0 0 0 0
1
0
0 0 13024 90
4 4511
-14 -60 14 -52
3 U15
38 -20 59 -12
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3417 0 0
2
5.89785e-315 5.43192e-315
0
4 4511
219 1037 241 0 20 29
0 26 27 28 29 2 62 62 67 66
65 64 68 69 70 0 0 0 0 0
5
0
0 0 13024 90
4 4511
-14 -60 14 -52
3 U16
38 -20 59 -12
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6882 0 0
2
5.89785e-315 5.43451e-315
0
7 Ground~
168 977 108 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7323 0 0
2
5.89785e-315 5.4371e-315
0
2 +V
167 945 292 0 1 3
0 63
0
0 0 54240 180
2 5V
7 -2 21 6
2 V6
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5262 0 0
2
5.89785e-315 5.43969e-315
0
7 Ground~
168 932 312 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7297 0 0
2
5.89785e-315 5.44228e-315
0
7 Ground~
168 1052 318 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
2
5.89785e-315 5.44487e-315
0
2 +V
167 1060 297 0 1 3
0 62
0
0 0 54240 180
2 5V
7 -2 21 6
2 V7
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7772 0 0
2
5.89785e-315 5.44746e-315
0
7 Ground~
168 536 102 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6238 0 0
2
42755.5 36
0
9 Inverter~
13 546 559 0 2 22
0 94 96
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U4E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
9459 0 0
2
42755.5 37
0
9 Inverter~
13 578 557 0 2 22
0 94 95
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U4D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3146 0 0
2
42755.5 38
0
9 Inverter~
13 514 555 0 2 22
0 94 97
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U4C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3236 0 0
2
42755.5 39
0
9 Inverter~
13 482 557 0 2 22
0 94 98
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U4B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3766 0 0
2
42755.5 40
0
7 Ground~
168 172 558 0 1 3
0 2
0
0 0 53344 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3921 0 0
2
42755.5 41
0
2 +V
167 170 535 0 1 3
0 99
0
0 0 54240 90
2 5V
-7 -15 7 -7
2 V5
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5622 0 0
2
42755.5 42
0
7 Ground~
168 204 485 0 1 3
0 2
0
0 0 53344 270
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
42755.5 43
0
9 2-In AND~
219 445 519 0 3 22
0 78 94 83
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
8101 0 0
2
42755.5 44
0
9 2-In AND~
219 349 518 0 3 22
0 81 94 93
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U12A
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7390 0 0
2
42755.5 45
0
9 2-In AND~
219 381 518 0 3 22
0 80 94 87
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5656 0 0
2
42755.5 46
0
9 2-In AND~
219 413 519 0 3 22
0 79 94 85
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6501 0 0
2
42755.5 47
0
9 2-In AND~
219 541 520 0 3 22
0 51 96 84
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U12C
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9939 0 0
2
42755.5 48
0
9 2-In AND~
219 509 519 0 3 22
0 52 97 86
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U12D
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
7700 0 0
2
42755.5 49
0
9 2-In AND~
219 477 519 0 3 22
0 11 98 88
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U13A
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
5463 0 0
2
42755.5 50
0
9 2-In AND~
219 573 520 0 3 22
0 50 95 82
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U12B
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
8614 0 0
2
42755.5 51
0
8 2-In OR~
219 394 458 0 3 22
0 93 88 89
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U11A
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3153 0 0
2
42755.5 52
0
8 2-In OR~
219 429 459 0 3 22
0 87 86 90
0
0 0 608 90
6 74LS32
-21 -24 21 -16
3 U9D
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
7372 0 0
2
42755.5 53
0
8 2-In OR~
219 462 460 0 3 22
0 85 84 91
0
0 0 608 90
6 74LS32
-21 -24 21 -16
3 U9C
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3974 0 0
2
42755.5 54
0
8 2-In OR~
219 497 461 0 3 22
0 83 82 92
0
0 0 608 90
6 74LS32
-21 -24 21 -16
3 U9B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4458 0 0
2
42755.5 55
0
4 4008
219 258 527 0 14 29
0 2 52 51 50 99 99 99 2 160
78 79 80 81 161
0
0 0 13024 0
4 4008
-14 -60 14 -52
3 U10
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
83 0 0
2
42755.5 56
0
7 Ground~
168 213 90 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6645 0 0
2
42755.5 57
0
8 2-In OR~
219 338 346 0 3 22
0 101 100 94
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3313 0 0
2
42755.5 58
0
9 2-In AND~
219 296 363 0 3 22
0 52 11 100
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3188 0 0
2
42755.5 59
0
9 2-In AND~
219 297 328 0 3 22
0 11 51 101
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3667 0 0
2
42755.5 60
0
4 4015
219 139 319 0 7 32
0 12 102 162 50 51 52 11
0
0 0 13024 0
4 4015
-14 -60 14 -52
3 U2A
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 5 4 3 10 7 9
6 5 4 3 10 15 1 14 13 12
11 2 0
65 0 0 512 2 1 1 0
1 U
8839 0 0
2
42755.5 61
0
9 2-In XOR~
219 207 201 0 3 22
0 51 103 10
0
0 0 608 180
6 74LS86
-21 -24 21 -16
3 U3A
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4966 0 0
2
42755.5 62
0
9 2-In XOR~
219 308 214 0 3 22
0 11 52 103
0
0 0 608 90
6 74LS86
-21 -24 21 -16
3 U3C
26 -3 47 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4293 0 0
2
42755.5 63
0
4 4511
219 311 130 0 20 29
0 2 2 2 94 2 111 111 110 109
108 107 106 105 104 0 0 0 0 0
1
0
0 0 13024 90
4 4511
-14 -60 14 -52
2 U6
41 -20 55 -12
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7459 0 0
2
42755.5 64
0
2 +V
167 371 167 0 1 3
0 111
0
0 0 54240 270
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7190 0 0
2
42755.5 65
0
7 Ground~
168 319 173 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
955 0 0
2
42755.5 66
0
9 CC 7-Seg~
183 490 136 0 17 19
10 104 105 106 107 108 109 110 163 2
0 1 1 0 0 0 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
493 0 0
2
42755.5 67
0
7 Ground~
168 501 397 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9550 0 0
2
42755.5 68
0
2 +V
167 536 377 0 1 3
0 121
0
0 0 54240 270
2 5V
-7 -15 7 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3398 0 0
2
42755.5 69
0
7 Pulser~
4 112 459 0 10 12
0 164 165 112 166 0 1 99 66 22
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5108 0 0
2
42755.5 70
0
4 4511
219 481 339 0 14 29
0 89 90 91 92 2 121 121 115 114
116 117 118 119 120
0
0 0 13024 90
4 4511
-14 -60 14 -52
2 U1
41 -20 55 -12
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7936 0 0
2
42755.5 71
0
9 CC 7-Seg~
183 580 138 0 17 19
10 120 119 118 117 116 114 115 167 2
1 1 1 1 1 1 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9993 0 0
2
42755.5 72
0
9 2-In AND~
219 162 396 0 3 22
0 113 112 102
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6682 0 0
2
42755.5 73
0
210
2 1 3 0 0 4224 0 2 52 0 0 2
786 315
786 283
0 1 4 0 0 4096 0 0 2 6 0 3
791 479
791 351
786 351
3 1 5 0 0 4224 0 4 51 0 0 4
833 391
833 261
809 261
809 253
2 2 6 0 0 4224 0 3 4 0 0 2
842 468
842 436
1 0 7 0 0 4096 0 3 0 0 8 2
842 504
861 504
0 1 4 0 0 0 0 0 4 9 0 3
734 479
824 479
824 436
3 1 8 0 0 4224 0 5 50 0 0 5
743 412
743 279
758 279
758 253
755 253
2 13 7 0 0 8320 0 5 49 0 0 4
752 457
861 457
861 664
851 664
1 15 4 0 0 4224 0 5 46 0 0 2
734 457
734 678
1 3 9 0 0 4224 0 7 6 0 0 2
78 198
100 198
2 3 10 0 0 4224 0 6 90 0 0 5
149 189
179 189
179 197
180 197
180 201
0 1 11 0 0 4096 0 0 6 187 0 5
181 283
181 213
154 213
154 207
149 207
2 1 12 0 0 4224 0 7 89 0 0 3
42 198
42 283
107 283
0 1 13 0 0 8320 0 0 38 30 0 5
1537 148
1537 217
1162 217
1162 264
1169 264
0 1 14 0 0 8320 0 0 37 31 0 5
1437 148
1437 222
1247 222
1247 263
1253 263
0 1 15 0 0 4224 0 0 36 32 0 3
1337 148
1337 263
1347 263
7 1 16 0 0 12416 0 44 35 0 0 5
1217 148
1231 148
1231 247
1433 247
1433 263
0 3 17 0 0 4224 0 0 41 19 0 4
1351 93
1463 93
1463 157
1471 157
0 3 17 0 0 0 0 0 42 20 0 4
1255 76
1351 76
1351 157
1376 157
0 3 17 0 0 0 0 0 43 21 0 4
1151 76
1255 76
1255 157
1277 157
3 3 17 0 0 0 0 39 44 0 0 4
1108 76
1151 76
1151 157
1169 157
0 4 18 0 0 4096 0 0 43 23 0 3
1269 148
1269 166
1277 166
3 2 18 0 0 4224 0 10 43 0 0 4
1364 72
1269 72
1269 148
1277 148
0 4 13 0 0 0 0 0 42 25 0 3
1364 148
1364 166
1376 166
0 2 13 0 0 0 0 0 42 30 0 4
1538 115
1364 115
1364 148
1376 148
4 0 19 0 0 4096 0 41 0 0 27 2
1471 166
1454 166
1 2 19 0 0 4224 0 8 41 0 0 3
1454 196
1454 148
1471 148
1 0 14 0 0 0 0 10 0 0 31 2
1409 81
1441 81
2 0 13 0 0 0 0 10 0 0 30 2
1409 63
1538 63
7 3 13 0 0 0 0 41 9 0 0 4
1519 148
1538 148
1538 37
1256 37
7 2 14 0 0 0 0 42 9 0 0 4
1424 148
1441 148
1441 46
1256 46
7 1 15 0 0 0 0 43 9 0 0 6
1325 148
1337 148
1337 91
1264 91
1264 55
1256 55
0 2 20 0 0 8192 0 0 44 34 0 3
1162 147
1162 148
1169 148
4 4 20 0 0 8320 0 9 44 0 0 4
1211 46
1162 46
1162 166
1169 166
0 9 21 0 0 12288 0 0 46 46 0 6
1216 650
1059 650
1059 774
646 774
646 714
664 714
0 10 22 0 0 8320 0 0 46 43 0 5
1051 640
1051 766
653 766
653 723
664 723
11 0 23 0 0 12416 0 46 0 0 44 5
664 732
659 732
659 759
1044 759
1044 631
0 12 24 0 0 8320 0 0 46 45 0 4
1037 621
1037 753
664 753
664 741
0 2 23 0 0 0 0 0 32 48 0 5
1370 434
1047 434
1047 473
977 473
977 457
0 2 22 0 0 0 0 0 31 47 0 5
1409 428
1041 428
1041 480
941 480
941 456
0 1 21 0 0 0 0 0 32 42 0 3
960 485
959 485
959 457
0 1 21 0 0 4224 0 0 31 46 0 5
1493 421
1035 421
1035 485
923 485
923 456
0 2 22 0 0 0 0 0 30 47 0 4
1246 640
946 640
946 537
973 537
3 0 23 0 0 0 0 30 0 0 48 4
973 546
950 546
950 631
1278 631
0 4 24 0 0 0 0 0 30 49 0 4
1311 621
960 621
960 555
973 555
4 1 21 0 0 0 0 35 24 0 0 5
1481 263
1493 263
1493 650
1214 650
1214 577
4 1 22 0 0 0 0 36 23 0 0 5
1395 263
1409 263
1409 640
1246 640
1246 577
1 4 23 0 0 0 0 22 37 0 0 7
1278 578
1278 631
1370 631
1370 347
1316 347
1316 263
1301 263
4 1 24 0 0 0 0 38 25 0 0 7
1217 264
1227 264
1227 354
1361 354
1361 621
1310 621
1310 578
2 0 25 0 0 4096 0 18 0 0 57 2
1200 577
1200 666
2 0 25 0 0 0 0 21 0 0 57 2
1168 577
1168 666
2 0 25 0 0 4096 0 20 0 0 57 2
1136 576
1136 666
2 0 25 0 0 0 0 19 0 0 57 2
1104 576
1104 666
1 0 25 0 0 0 0 14 0 0 57 2
1232 612
1232 666
1 0 25 0 0 0 0 13 0 0 57 2
1264 610
1264 666
1 0 25 0 0 0 0 11 0 0 57 2
1296 614
1296 666
3 1 25 0 0 20624 0 33 12 0 0 7
950 350
994 350
994 464
1069 464
1069 666
1328 666
1328 612
3 4 25 0 0 0 0 33 57 0 0 3
950 350
921 350
921 258
3 1 26 0 0 8320 0 26 58 0 0 4
1144 465
1144 384
1010 384
1010 258
2 3 27 0 0 8320 0 58 27 0 0 4
1019 258
1019 380
1179 380
1179 466
3 3 28 0 0 8320 0 28 58 0 0 4
1212 467
1212 374
1028 374
1028 258
4 3 29 0 0 8320 0 58 29 0 0 4
1037 258
1037 370
1247 370
1247 468
10 1 30 0 0 12416 0 30 18 0 0 5
1037 573
1046 573
1046 609
1182 609
1182 577
11 1 31 0 0 12416 0 30 21 0 0 5
1037 564
1051 564
1051 601
1150 601
1150 577
1 12 32 0 0 8320 0 20 30 0 0 5
1118 576
1118 584
1056 584
1056 555
1037 555
13 1 33 0 0 8320 0 30 19 0 0 4
1037 546
1060 546
1060 576
1086 576
2 3 34 0 0 4224 0 29 25 0 0 3
1256 514
1319 514
1319 533
3 1 35 0 0 12416 0 18 29 0 0 4
1191 532
1213 532
1213 514
1238 514
3 2 36 0 0 8320 0 22 28 0 0 4
1287 533
1287 520
1221 520
1221 513
3 1 37 0 0 8320 0 21 28 0 0 4
1159 532
1159 519
1203 519
1203 513
3 2 38 0 0 8320 0 23 27 0 0 4
1255 532
1255 524
1188 524
1188 512
3 1 39 0 0 8320 0 20 27 0 0 4
1127 531
1127 515
1170 515
1170 512
3 2 40 0 0 8320 0 24 26 0 0 4
1223 532
1223 528
1153 528
1153 511
3 1 41 0 0 8320 0 19 26 0 0 3
1095 531
1095 511
1135 511
2 2 42 0 0 4224 0 12 25 0 0 2
1328 576
1328 578
2 2 43 0 0 0 0 11 22 0 0 2
1296 578
1296 578
2 2 44 0 0 4224 0 13 23 0 0 2
1264 574
1264 577
2 2 45 0 0 4224 0 14 24 0 0 2
1232 576
1232 577
1 8 2 0 0 4096 0 15 30 0 0 4
926 596
954 596
954 591
973 591
0 7 46 0 0 16384 0 0 30 81 0 5
964 573
964 578
965 578
965 582
973 582
0 6 46 0 0 8192 0 0 30 82 0 3
964 570
964 573
973 573
1 5 46 0 0 4224 0 16 30 0 0 4
928 570
965 570
965 564
973 564
1 1 2 0 0 0 0 17 30 0 0 4
958 523
965 523
965 528
973 528
3 2 47 0 0 4224 0 32 33 0 0 3
968 412
968 396
959 396
3 1 48 0 0 4224 0 31 33 0 0 3
932 411
932 396
941 396
2 0 49 0 0 8192 0 35 0 0 89 3
1433 281
1417 281
1417 227
2 0 49 0 0 0 0 36 0 0 89 3
1347 281
1325 281
1325 227
0 2 49 0 0 0 0 0 37 89 0 3
1235 227
1235 281
1253 281
3 2 49 0 0 12416 0 34 38 0 0 6
1534 259
1512 259
1512 227
1156 227
1156 282
1169 282
0 8 50 0 0 8192 0 0 46 134 0 3
433 603
433 705
664 705
0 7 51 0 0 8192 0 0 46 135 0 3
442 597
442 696
664 696
0 6 52 0 0 8192 0 0 46 136 0 3
452 592
452 687
664 687
0 5 11 0 0 8192 0 0 46 137 0 3
461 588
461 678
664 678
0 3 2 0 0 0 0 0 46 95 0 3
663 651
663 660
670 660
1 2 2 0 0 0 0 48 46 0 0 3
663 635
663 651
670 651
0 4 53 0 0 4224 0 0 46 98 0 3
647 642
647 669
670 669
14 1 2 0 0 0 0 46 45 0 0 3
734 651
734 648
747 648
1 1 53 0 0 0 0 46 47 0 0 3
670 642
647 642
647 636
1 4 54 0 0 12416 0 49 54 0 0 4
787 610
787 563
681 563
681 265
3 2 55 0 0 4224 0 54 49 0 0 5
675 265
675 572
767 572
767 619
787 619
3 2 56 0 0 16512 0 49 54 0 0 5
787 628
759 628
759 580
669 580
669 265
1 4 57 0 0 4224 0 54 49 0 0 5
663 265
663 586
754 586
754 637
787 637
22 8 58 0 0 8320 0 46 49 0 0 3
740 741
787 741
787 673
7 21 59 0 0 8320 0 49 46 0 0 4
787 664
781 664
781 732
740 732
20 6 60 0 0 8320 0 46 49 0 0 4
740 723
776 723
776 655
787 655
19 5 61 0 0 8320 0 46 49 0 0 4
740 714
773 714
773 646
787 646
0 2 2 0 0 0 0 0 51 108 0 3
786 225
809 225
809 233
2 0 2 0 0 0 0 50 0 0 109 3
755 233
755 225
783 225
2 1 2 0 0 8192 0 52 53 0 0 3
786 263
783 263
783 212
0 1 62 0 0 4224 0 0 63 111 0 2
1060 273
1060 282
6 7 62 0 0 0 0 58 58 0 0 4
1055 264
1055 273
1064 273
1064 264
1 5 2 0 0 0 0 62 58 0 0 4
1052 312
1052 294
1046 294
1046 264
1 5 2 0 0 0 0 61 57 0 0 3
932 306
930 306
930 264
6 0 63 0 0 4224 0 57 0 0 115 3
939 264
939 271
945 271
1 7 63 0 0 0 0 60 57 0 0 4
945 277
945 271
948 271
948 264
4 11 64 0 0 4224 0 56 58 0 0 4
1023 174
1023 188
1037 188
1037 194
5 10 65 0 0 16512 0 56 58 0 0 6
1029 174
1029 178
1031 178
1031 184
1046 184
1046 194
9 6 66 0 0 8320 0 58 56 0 0 4
1055 194
1055 181
1035 181
1035 174
7 8 67 0 0 8320 0 56 58 0 0 4
1041 174
1041 177
1064 177
1064 194
3 12 68 0 0 8320 0 56 58 0 0 4
1017 174
1017 183
1028 183
1028 194
2 13 69 0 0 4224 0 56 58 0 0 4
1011 174
1011 189
1019 189
1019 194
1 14 70 0 0 4224 0 56 58 0 0 3
1005 174
1005 194
1010 194
4 11 71 0 0 4224 0 55 57 0 0 3
925 173
925 194
921 194
3 12 72 0 0 4224 0 55 57 0 0 4
919 173
919 186
912 186
912 194
5 10 73 0 0 8320 0 55 57 0 0 3
931 173
930 173
930 194
6 9 74 0 0 12416 0 55 57 0 0 4
937 173
937 179
939 179
939 194
8 7 75 0 0 4224 0 57 55 0 0 4
948 194
948 176
943 176
943 173
13 2 76 0 0 4224 0 57 55 0 0 4
903 194
903 181
913 181
913 173
14 1 77 0 0 4224 0 57 55 0 0 4
894 194
894 176
907 176
907 173
0 1 2 0 0 0 0 0 59 131 0 3
979 96
977 96
977 102
9 9 2 0 0 8320 0 55 56 0 0 3
928 95
928 96
1026 96
1 9 2 0 0 0 0 64 100 0 0 2
536 96
580 96
9 1 2 0 0 0 0 95 64 0 0 3
490 94
490 96
536 96
0 1 50 0 0 20608 0 0 79 173 0 7
212 313
261 313
261 219
47 219
47 603
563 603
563 541
0 1 51 0 0 16512 0 0 76 178 0 6
219 337
219 227
54 227
54 597
531 597
531 541
0 1 52 0 0 16512 0 0 77 186 0 6
226 295
226 234
60 234
60 592
499 592
499 540
0 1 11 0 0 16512 0 0 78 187 0 6
235 286
235 242
68 242
68 588
467 588
467 540
10 1 78 0 0 12416 0 84 72 0 0 5
290 536
299 536
299 572
435 572
435 540
11 1 79 0 0 12416 0 84 75 0 0 5
290 527
304 527
304 564
403 564
403 540
1 12 80 0 0 8320 0 74 84 0 0 5
371 539
371 547
309 547
309 518
290 518
13 1 81 0 0 8320 0 84 73 0 0 4
290 509
313 509
313 539
339 539
2 3 82 0 0 4224 0 83 79 0 0 3
509 477
572 477
572 496
3 1 83 0 0 12416 0 72 83 0 0 4
444 495
466 495
466 477
491 477
3 2 84 0 0 8320 0 76 82 0 0 4
540 496
540 483
474 483
474 476
3 1 85 0 0 8320 0 75 82 0 0 4
412 495
412 482
456 482
456 476
3 2 86 0 0 8320 0 77 81 0 0 4
508 495
508 487
441 487
441 475
3 1 87 0 0 8320 0 74 81 0 0 4
380 494
380 478
423 478
423 475
3 2 88 0 0 8320 0 78 80 0 0 4
476 495
476 491
406 491
406 474
1 3 89 0 0 4224 0 99 80 0 0 4
454 356
454 414
397 414
397 428
3 2 90 0 0 12416 0 81 99 0 0 6
432 429
432 419
460 419
460 383
463 383
463 356
3 3 91 0 0 4224 0 99 82 0 0 4
472 356
472 422
465 422
465 430
3 4 92 0 0 12416 0 83 99 0 0 4
500 431
500 420
481 420
481 356
3 1 93 0 0 8320 0 73 80 0 0 3
348 494
348 474
388 474
1 0 94 0 0 4096 0 65 0 0 157 2
549 577
549 584
1 0 94 0 0 4096 0 68 0 0 157 2
485 575
485 584
1 0 94 0 0 4096 0 67 0 0 157 2
517 573
517 584
0 1 94 0 0 8192 0 0 66 165 0 4
452 553
452 584
581 584
581 575
2 2 95 0 0 4224 0 66 79 0 0 2
581 539
581 541
2 2 96 0 0 0 0 65 76 0 0 2
549 541
549 541
2 2 97 0 0 4224 0 67 77 0 0 2
517 537
517 540
2 2 98 0 0 4224 0 68 78 0 0 2
485 539
485 540
2 0 94 0 0 0 0 73 0 0 165 2
357 539
357 553
2 0 94 0 0 0 0 74 0 0 165 2
389 539
389 553
2 0 94 0 0 0 0 75 0 0 165 2
421 540
421 553
0 2 94 0 0 12416 0 0 72 177 0 6
383 344
383 406
319 406
319 553
453 553
453 540
1 8 2 0 0 0 0 69 84 0 0 4
179 559
207 559
207 554
226 554
0 7 99 0 0 16384 0 0 84 168 0 5
217 536
217 541
218 541
218 545
226 545
0 6 99 0 0 8192 0 0 84 169 0 3
217 533
217 536
226 536
1 5 99 0 0 4224 0 70 84 0 0 4
181 533
218 533
218 527
226 527
1 1 2 0 0 0 0 71 84 0 0 4
211 486
218 486
218 491
226 491
0 2 52 0 0 0 0 0 84 186 0 5
249 295
249 464
180 464
180 500
226 500
0 3 51 0 0 0 0 0 84 178 0 5
241 337
241 457
172 457
172 509
226 509
4 4 50 0 0 0 0 89 84 0 0 6
171 310
212 310
212 450
167 450
167 518
226 518
0 1 2 0 0 0 0 0 92 176 0 2
284 153
284 147
2 0 2 0 0 0 0 92 0 0 176 2
293 147
293 153
1 3 2 0 0 0 0 85 92 0 0 5
213 98
211 98
211 153
302 153
302 147
4 3 94 0 0 0 0 92 86 0 0 7
311 147
311 159
333 159
333 306
383 306
383 346
371 346
2 5 51 0 0 0 0 88 89 0 0 5
273 337
219 337
219 302
171 302
171 301
0 1 52 0 0 0 0 0 87 186 0 3
265 295
265 354
272 354
1 0 11 0 0 0 0 88 0 0 181 2
273 319
256 319
0 2 11 0 0 0 0 0 87 187 0 3
256 286
256 372
272 372
3 2 100 0 0 4224 0 87 86 0 0 3
317 363
317 355
325 355
3 1 101 0 0 4224 0 88 86 0 0 3
318 328
318 337
325 337
3 2 102 0 0 8320 0 101 89 0 0 5
183 396
183 340
90 340
90 292
107 292
5 1 51 0 0 0 0 89 90 0 0 4
171 301
241 301
241 210
229 210
2 6 52 0 0 0 0 91 89 0 0 5
320 233
320 295
226 295
226 292
171 292
7 1 11 0 0 0 0 89 91 0 0 5
171 283
205 283
205 286
302 286
302 233
2 3 103 0 0 4224 0 90 91 0 0 5
229 192
287 192
287 179
311 179
311 184
14 1 104 0 0 8320 0 92 95 0 0 6
284 83
284 55
424 55
424 171
469 171
469 172
2 13 105 0 0 16512 0 95 92 0 0 6
475 172
475 176
419 176
419 58
293 58
293 83
12 3 106 0 0 12416 0 92 95 0 0 6
302 83
302 61
412 61
412 180
481 180
481 172
4 11 107 0 0 12416 0 95 92 0 0 6
487 172
487 184
406 184
406 67
311 67
311 83
10 5 108 0 0 12416 0 92 95 0 0 6
320 83
320 72
399 72
399 187
493 187
493 172
6 9 109 0 0 12416 0 95 92 0 0 6
499 172
499 192
392 192
392 77
329 77
329 83
8 7 110 0 0 12416 0 92 95 0 0 5
338 83
386 83
386 196
505 196
505 172
5 1 2 0 0 0 0 92 94 0 0 4
320 153
320 159
319 159
319 167
0 6 111 0 0 8192 0 0 92 198 0 3
338 157
338 153
329 153
7 1 111 0 0 8320 0 92 93 0 0 5
338 153
338 157
352 157
352 166
359 166
3 2 112 0 0 4224 0 98 101 0 0 3
136 450
136 405
138 405
1 1 113 0 0 8320 0 1 101 0 0 4
124 377
130 377
130 387
138 387
6 9 114 0 0 4224 0 100 99 0 0 6
589 174
589 266
500 266
500 286
499 286
499 292
8 7 115 0 0 12416 0 99 100 0 0 4
508 292
508 274
595 274
595 174
10 5 116 0 0 8320 0 99 100 0 0 4
490 292
490 260
583 260
583 174
11 4 117 0 0 8320 0 99 100 0 0 4
481 292
481 251
577 251
577 174
12 3 118 0 0 8320 0 99 100 0 0 4
472 292
472 245
571 245
571 174
2 13 119 0 0 8320 0 100 99 0 0 4
565 174
565 235
463 235
463 292
14 1 120 0 0 8320 0 99 100 0 0 4
454 292
454 228
559 228
559 174
0 6 121 0 0 8192 0 0 99 210 0 3
508 376
499 376
499 362
1 5 2 0 0 0 0 96 99 0 0 3
501 391
490 391
490 362
1 7 121 0 0 4224 0 97 99 0 0 3
524 376
508 376
508 362
5
-27 0 0 0 400 0 0 0 0 0 0 0 49
11 Courier New
0 32768 0 3
674 587 723 616
674 587 723 616
3 ULA
-24 0 0 0 400 0 0 0 0 0 0 0 49
11 Courier New
0 0 0 4
93 91 162 129
102 95 157 121
4 LFSR
-24 0 0 0 400 0 0 0 0 0 0 0 49
11 Courier New
0 0 0 11
451 37 616 107
464 40 615 92
11 1o Operando
-24 0 0 0 400 0 0 0 0 0 0 0 49
11 Courier New
0 0 0 11
893 43 1058 81
905 47 1056 73
11 2o Operando
-27 0 0 0 400 0 0 0 0 0 0 0 49
11 Courier New
0 32768 0 11
647 152 820 181
647 152 820 181
11 INTERATIVOS
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1573236 1472576 100 100 0 0
0 0 0 0
65 211 226 281
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 5e-17
1
300 145
0 2 0 0 3	0 211 0 0
5112028 8550976 100 100 0 0
77 66 1277 246
65 419 1366 752
1277 66
77 66
1277 66
1277 246
0 0
0 0 0 0 0 0
12409 0
4 1 200
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
